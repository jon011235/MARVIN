/*
    Project:    MARVIN
    Sector:     CPU
    Summary:    Central processing unit, consisting of cu and alu
    Authors:    Leonard Pfeiffer
*/

module cpu(
    input clk
);

endmodule