/*
    Project:    MARVIN
    Sector:     CPU
    Summary:    Control unit, manager for interactions between other
    Authors:    Leonard Pfeiffer
*/

module cu(
    input clk
);

endmodule