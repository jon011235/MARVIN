/*
    Project:    MARVIN
    Sector:     CPU
    Summary:    Types and constants for the cpu
    Authors:    Leonard Pfeiffer
*/

package cpu_pkg

endpackage