/*
    Project:    MARVIN
    Sector:     CPU
    Summary:    Arithmetical logic unit, for calculations
    Authors:    Leonard Pfeiffer
*/

module alu(
    input clk
);

endmodule