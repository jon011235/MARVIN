/*
    Project:    MARVIN
    Sector:     COM
    Summary:    Uart interface package
    Authors:    Leonard Pfeiffer
*/

package uart_pkg;
    typedef enum {NONE, EVEN, ODD, MARK, SPACE} parity_t;
endpackage